
endmodule: noc

endpackage: noc