package noc;

import toplevel_defs::*;

import chain_l2::*;
import ring_l2::*;
import mesh_l2::*;
import folrus_l2::*;
//import butterfly_l2::*;
import hypercube_l2::*;

module noc (Empty);
